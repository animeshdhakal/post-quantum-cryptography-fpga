package ntt_rom_pkg;
    // Zetas in Montgomery Domain (x * 2^16 mod 3329)
    // Order matches Cooley-Tukey processing order (k=1..127)
    function automatic logic [15:0] get_zeta(input logic [6:0] idx);
        case (idx)
            7'd0: return 16'd2285;
            7'd1: return 16'd2571;
            7'd2: return 16'd2970;
            7'd3: return 16'd1812;
            7'd4: return 16'd1493;
            7'd5: return 16'd1422;
            7'd6: return 16'd287;
            7'd7: return 16'd202;
            7'd8: return 16'd3158;
            7'd9: return 16'd622;
            7'd10: return 16'd1577;
            7'd11: return 16'd182;
            7'd12: return 16'd962;
            7'd13: return 16'd2127;
            7'd14: return 16'd1855;
            7'd15: return 16'd1468;
            7'd16: return 16'd573;
            7'd17: return 16'd2004;
            7'd18: return 16'd264;
            7'd19: return 16'd383;
            7'd20: return 16'd2500;
            7'd21: return 16'd1458;
            7'd22: return 16'd1727;
            7'd23: return 16'd3199;
            7'd24: return 16'd2648;
            7'd25: return 16'd1017;
            7'd26: return 16'd732;
            7'd27: return 16'd608;
            7'd28: return 16'd1787;
            7'd29: return 16'd411;
            7'd30: return 16'd3124;
            7'd31: return 16'd1758;
            7'd32: return 16'd1223;
            7'd33: return 16'd652;
            7'd34: return 16'd2777;
            7'd35: return 16'd1015;
            7'd36: return 16'd2036;
            7'd37: return 16'd1491;
            7'd38: return 16'd3047;
            7'd39: return 16'd1785;
            7'd40: return 16'd516;
            7'd41: return 16'd3321;
            7'd42: return 16'd3009;
            7'd43: return 16'd2663;
            7'd44: return 16'd1711;
            7'd45: return 16'd2167;
            7'd46: return 16'd126;
            7'd47: return 16'd1469;
            7'd48: return 16'd2476;
            7'd49: return 16'd3239;
            7'd50: return 16'd3058;
            7'd51: return 16'd830;
            7'd52: return 16'd107;
            7'd53: return 16'd1908;
            7'd54: return 16'd3082;
            7'd55: return 16'd2378;
            7'd56: return 16'd2931;
            7'd57: return 16'd961;
            7'd58: return 16'd1821;
            7'd59: return 16'd2604;
            7'd60: return 16'd448;
            7'd61: return 16'd2264;
            7'd62: return 16'd677;
            7'd63: return 16'd2054;
            7'd64: return 16'd2226;
            7'd65: return 16'd430;
            7'd66: return 16'd555;
            7'd67: return 16'd843;
            7'd68: return 16'd2078;
            7'd69: return 16'd871;
            7'd70: return 16'd1550;
            7'd71: return 16'd105;
            7'd72: return 16'd422;
            7'd73: return 16'd587;
            7'd74: return 16'd177;
            7'd75: return 16'd3094;
            7'd76: return 16'd3038;
            7'd77: return 16'd2869;
            7'd78: return 16'd1574;
            7'd79: return 16'd1653;
            7'd80: return 16'd3083;
            7'd81: return 16'd778;
            7'd82: return 16'd1159;
            7'd83: return 16'd3182;
            7'd84: return 16'd2552;
            7'd85: return 16'd1483;
            7'd86: return 16'd2727;
            7'd87: return 16'd1119;
            7'd88: return 16'd1739;
            7'd89: return 16'd644;
            7'd90: return 16'd2457;
            7'd91: return 16'd349;
            7'd92: return 16'd418;
            7'd93: return 16'd329;
            7'd94: return 16'd3173;
            7'd95: return 16'd3254;
            7'd96: return 16'd817;
            7'd97: return 16'd1097;
            7'd98: return 16'd603;
            7'd99: return 16'd610;
            7'd100: return 16'd1322;
            7'd101: return 16'd2044;
            7'd102: return 16'd1864;
            7'd103: return 16'd384;
            7'd104: return 16'd2114;
            7'd105: return 16'd3193;
            7'd106: return 16'd1218;
            7'd107: return 16'd1994;
            7'd108: return 16'd2455;
            7'd109: return 16'd220;
            7'd110: return 16'd2142;
            7'd111: return 16'd1670;
            7'd112: return 16'd2144;
            7'd113: return 16'd1799;
            7'd114: return 16'd2051;
            7'd115: return 16'd794;
            7'd116: return 16'd1819;
            7'd117: return 16'd2475;
            7'd118: return 16'd2459;
            7'd119: return 16'd478;
            7'd120: return 16'd3221;
            7'd121: return 16'd3021;
            7'd122: return 16'd996;
            7'd123: return 16'd991;
            7'd124: return 16'd958;
            7'd125: return 16'd1869;
            7'd126: return 16'd1522;
            7'd127: return 16'd1628;
            default: return 16'd0;
        endcase
    endfunction
endpackage
